///////////////////////////////////////////
// cdc_sync_stb.sv
//
// Written: james.stine@okstate.edu, jacob.pease@okstate.edu, matotto@okstate.edu 28 July 2025
// Modified: 
//
// Purpose: CDC synchronizer
// 
// A component of the CORE-V-WALLY configurable RISC-V project.
// https://github.com/openhwgroup/cvw
// 
// Copyright (C) 2021-25 Harvey Mudd College & Oklahoma State University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

module cdc_sync_stb #(parameter RISING_EDGE = 1)
   (input logic  a,
    input logic  clk_b,
    output logic b);

   logic 	 sync1, sync2;
   logic 	 lock;
   
   initial
     lock = 0;
   
   always @(posedge clk_b) begin
      sync1 <= a;
      sync2 <= sync1;
      
      if (RISING_EDGE) begin
         if (sync2 && ~lock) begin
            lock <= 1;
            b <= 1;
         end
         if (b)
           b <= 0;
         if (~sync2)
           lock <= 0;
      end else begin
         if (~sync2 && ~lock) begin
            lock <= 1;
            b <= 0;
         end
         if (~b)
           b <= 1;
         if (sync2)
           lock <= 0;
      end
   end
   
endmodule // cdc_sync_stb

